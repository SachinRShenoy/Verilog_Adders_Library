`ifndef PARAMS_VH
`define PARAMS_VH

`define N 8

`endif
